LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.CONSTANTS.ALL;
USE WORK.LIBNODE.ALL;


ENTITY NoC IS
	PORT (SW			: IN STD_LOGIC_VECTOR(17 DOWNTO 0);
			CLOCK_50	: IN STD_LOGIC;
			LEDR		: OUT STD_LOGIC_VECTOR(17 DOWNTO 0));
END;

ARCHITECTURE STRUCTURE OF NoC IS

component NOCUNIT
generic (id : integer; count : integer; nocdim : STD_LOGIC_VECTOR(63 downto 0));
PORT (	Clk 					: IN std_logic;
	rst_n 					: IN std_logic;				
	NorthOut				: OUT P_PORT_VERTICAL;
	SouthIn				: IN  P_PORT_VERTICAL;
	EastOut	   		: OUT P_PORT_HORIZONTAL;
	WestIn				: IN  P_PORT_HORIZONTAL;							
	CoreAddress			: IN  Address					
	);
END component;



-------------------------------------------------
--SIGNALS for NODE 000000

SIGNAL N_000000EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_000000NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_000000CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 000001

SIGNAL N_000001EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_000001NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_000001CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 000010

SIGNAL N_000010EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_000010NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_000010CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 000011

SIGNAL N_000011EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_000011NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_000011CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 000100

SIGNAL N_000100EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_000100NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_000100CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 001000

SIGNAL N_001000EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_001000NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_001000CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 001001

SIGNAL N_001001EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_001001NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_001001CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 001010

SIGNAL N_001010EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_001010NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_001010CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 001011

SIGNAL N_001011EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_001011NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_001011CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 001100

SIGNAL N_001100EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_001100NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_001100CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 010000

SIGNAL N_010000EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_010000NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_010000CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 010001

SIGNAL N_010001EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_010001NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_010001CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 010010

SIGNAL N_010010EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_010010NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_010010CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 010011

SIGNAL N_010011EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_010011NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_010011CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 010100

SIGNAL N_010100EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_010100NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_010100CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 011000

SIGNAL N_011000EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_011000NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_011000CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 011001

SIGNAL N_011001EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_011001NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_011001CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 011010

SIGNAL N_011010EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_011010NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_011010CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 011011

SIGNAL N_011011EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_011011NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_011011CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 011100

SIGNAL N_011100EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_011100NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_011100CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 100000

SIGNAL N_100000EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_100000NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_100000CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 100001

SIGNAL N_100001EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_100001NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_100001CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 100010

SIGNAL N_100010EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_100010NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_100010CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 100011

SIGNAL N_100011EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_100011NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_100011CORE_ADDRESS			:Address;

-------------------------------------------------
--SIGNALS for NODE 100100

SIGNAL N_100100EAST_OUT			:P_PORT_HORIZONTAL;
SIGNAL N_100100NORTH_OUT			:P_PORT_VERTICAL;
SIGNAL N_100100CORE_ADDRESS			:Address;




begin
	NOCUNIT000000 : NOCUNIT
generic map ( id => 0, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_000000NORTH_OUT,
				N_000001NORTH_OUT,
				N_000000EAST_OUT,
				N_100000EAST_OUT,
				N_000000CORE_ADDRESS);
	NOCUNIT000001 : NOCUNIT
generic map ( id => 5, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_000001NORTH_OUT,
				N_000010NORTH_OUT,
				N_000001EAST_OUT,
				N_100001EAST_OUT,
				N_000001CORE_ADDRESS);
	NOCUNIT000010 : NOCUNIT
generic map ( id => 10, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_000010NORTH_OUT,
				N_000011NORTH_OUT,
				N_000010EAST_OUT,
				N_100010EAST_OUT,
				N_000010CORE_ADDRESS);
	NOCUNIT000011 : NOCUNIT
generic map ( id => 15, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_000011NORTH_OUT,
				N_000100NORTH_OUT,
				N_000011EAST_OUT,
				N_100011EAST_OUT,
				N_000011CORE_ADDRESS);
	NOCUNIT000100 : NOCUNIT
generic map ( id => 20, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_000100NORTH_OUT,
				N_000000NORTH_OUT,
				N_000100EAST_OUT,
				N_100100EAST_OUT,
				N_000100CORE_ADDRESS);
	NOCUNIT001000 : NOCUNIT
generic map ( id => 1, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_001000NORTH_OUT,
				N_001001NORTH_OUT,
				N_001000EAST_OUT,
				N_000000EAST_OUT,
				N_001000CORE_ADDRESS);
	NOCUNIT001001 : NOCUNIT
generic map ( id => 6, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_001001NORTH_OUT,
				N_001010NORTH_OUT,
				N_001001EAST_OUT,
				N_000001EAST_OUT,
				N_001001CORE_ADDRESS);
	NOCUNIT001010 : NOCUNIT
generic map ( id => 11, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_001010NORTH_OUT,
				N_001011NORTH_OUT,
				N_001010EAST_OUT,
				N_000010EAST_OUT,
				N_001010CORE_ADDRESS);
	NOCUNIT001011 : NOCUNIT
generic map ( id => 16, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_001011NORTH_OUT,
				N_001100NORTH_OUT,
				N_001011EAST_OUT,
				N_000011EAST_OUT,
				N_001011CORE_ADDRESS);
	NOCUNIT001100 : NOCUNIT
generic map ( id => 21, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_001100NORTH_OUT,
				N_001000NORTH_OUT,
				N_001100EAST_OUT,
				N_000100EAST_OUT,
				N_001100CORE_ADDRESS);
	NOCUNIT010000 : NOCUNIT
generic map ( id => 2, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_010000NORTH_OUT,
				N_010001NORTH_OUT,
				N_010000EAST_OUT,
				N_001000EAST_OUT,
				N_010000CORE_ADDRESS);
	NOCUNIT010001 : NOCUNIT
generic map ( id => 7, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_010001NORTH_OUT,
				N_010010NORTH_OUT,
				N_010001EAST_OUT,
				N_001001EAST_OUT,
				N_010001CORE_ADDRESS);
	NOCUNIT010010 : NOCUNIT
generic map ( id => 12, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_010010NORTH_OUT,
				N_010011NORTH_OUT,
				N_010010EAST_OUT,
				N_001010EAST_OUT,
				N_010010CORE_ADDRESS);
	NOCUNIT010011 : NOCUNIT
generic map ( id => 17, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_010011NORTH_OUT,
				N_010100NORTH_OUT,
				N_010011EAST_OUT,
				N_001011EAST_OUT,
				N_010011CORE_ADDRESS);
	NOCUNIT010100 : NOCUNIT
generic map ( id => 22, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_010100NORTH_OUT,
				N_010000NORTH_OUT,
				N_010100EAST_OUT,
				N_001100EAST_OUT,
				N_010100CORE_ADDRESS);
	NOCUNIT011000 : NOCUNIT
generic map ( id => 3, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_011000NORTH_OUT,
				N_011001NORTH_OUT,
				N_011000EAST_OUT,
				N_010000EAST_OUT,
				N_011000CORE_ADDRESS);
	NOCUNIT011001 : NOCUNIT
generic map ( id => 8, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_011001NORTH_OUT,
				N_011010NORTH_OUT,
				N_011001EAST_OUT,
				N_010001EAST_OUT,
				N_011001CORE_ADDRESS);
	NOCUNIT011010 : NOCUNIT
generic map ( id => 13, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_011010NORTH_OUT,
				N_011011NORTH_OUT,
				N_011010EAST_OUT,
				N_010010EAST_OUT,
				N_011010CORE_ADDRESS);
	NOCUNIT011011 : NOCUNIT
generic map ( id => 18, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_011011NORTH_OUT,
				N_011100NORTH_OUT,
				N_011011EAST_OUT,
				N_010011EAST_OUT,
				N_011011CORE_ADDRESS);
	NOCUNIT011100 : NOCUNIT
generic map ( id => 23, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_011100NORTH_OUT,
				N_011000NORTH_OUT,
				N_011100EAST_OUT,
				N_010100EAST_OUT,
				N_011100CORE_ADDRESS);
	NOCUNIT100000 : NOCUNIT
generic map ( id => 4, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_100000NORTH_OUT,
				N_100001NORTH_OUT,
				N_100000EAST_OUT,
				N_011000EAST_OUT,
				N_100000CORE_ADDRESS);
	NOCUNIT100001 : NOCUNIT
generic map ( id => 9, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_100001NORTH_OUT,
				N_100010NORTH_OUT,
				N_100001EAST_OUT,
				N_011001EAST_OUT,
				N_100001CORE_ADDRESS);
	NOCUNIT100010 : NOCUNIT
generic map ( id => 14, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_100010NORTH_OUT,
				N_100011NORTH_OUT,
				N_100010EAST_OUT,
				N_011010EAST_OUT,
				N_100010CORE_ADDRESS);
	NOCUNIT100011 : NOCUNIT
generic map ( id => 19, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_100011NORTH_OUT,
				N_100100NORTH_OUT,
				N_100011EAST_OUT,
				N_011011EAST_OUT,
				N_100011CORE_ADDRESS);
	NOCUNIT100100 : NOCUNIT
generic map ( id => 24, count => 25, nocdim => x"0001000100050005" )
 port map( 
				CLOCK_50,
				SW(17),
				N_100100NORTH_OUT,
				N_100000NORTH_OUT,
				N_100100EAST_OUT,
				N_011100EAST_OUT,
				N_100100CORE_ADDRESS);








	N_000000CORE_ADDRESS.X <= "000";
	N_000000CORE_ADDRESS.Y <= "000";
	N_000001CORE_ADDRESS.X <= "000";
	N_000001CORE_ADDRESS.Y <= "001";
	N_000010CORE_ADDRESS.X <= "000";
	N_000010CORE_ADDRESS.Y <= "010";
	N_000011CORE_ADDRESS.X <= "000";
	N_000011CORE_ADDRESS.Y <= "011";
	N_000100CORE_ADDRESS.X <= "000";
	N_000100CORE_ADDRESS.Y <= "100";
	N_001000CORE_ADDRESS.X <= "001";
	N_001000CORE_ADDRESS.Y <= "000";
	N_001001CORE_ADDRESS.X <= "001";
	N_001001CORE_ADDRESS.Y <= "001";
	N_001010CORE_ADDRESS.X <= "001";
	N_001010CORE_ADDRESS.Y <= "010";
	N_001011CORE_ADDRESS.X <= "001";
	N_001011CORE_ADDRESS.Y <= "011";
	N_001100CORE_ADDRESS.X <= "001";
	N_001100CORE_ADDRESS.Y <= "100";
	N_010000CORE_ADDRESS.X <= "010";
	N_010000CORE_ADDRESS.Y <= "000";
	N_010001CORE_ADDRESS.X <= "010";
	N_010001CORE_ADDRESS.Y <= "001";
	N_010010CORE_ADDRESS.X <= "010";
	N_010010CORE_ADDRESS.Y <= "010";
	N_010011CORE_ADDRESS.X <= "010";
	N_010011CORE_ADDRESS.Y <= "011";
	N_010100CORE_ADDRESS.X <= "010";
	N_010100CORE_ADDRESS.Y <= "100";
	N_011000CORE_ADDRESS.X <= "011";
	N_011000CORE_ADDRESS.Y <= "000";
	N_011001CORE_ADDRESS.X <= "011";
	N_011001CORE_ADDRESS.Y <= "001";
	N_011010CORE_ADDRESS.X <= "011";
	N_011010CORE_ADDRESS.Y <= "010";
	N_011011CORE_ADDRESS.X <= "011";
	N_011011CORE_ADDRESS.Y <= "011";
	N_011100CORE_ADDRESS.X <= "011";
	N_011100CORE_ADDRESS.Y <= "100";
	N_100000CORE_ADDRESS.X <= "100";
	N_100000CORE_ADDRESS.Y <= "000";
	N_100001CORE_ADDRESS.X <= "100";
	N_100001CORE_ADDRESS.Y <= "001";
	N_100010CORE_ADDRESS.X <= "100";
	N_100010CORE_ADDRESS.Y <= "010";
	N_100011CORE_ADDRESS.X <= "100";
	N_100011CORE_ADDRESS.Y <= "011";
	N_100100CORE_ADDRESS.X <= "100";
	N_100100CORE_ADDRESS.Y <= "100";
end; 

