LIBRARY ieee;
USE ieee.std_logic_1164.all; 
use work.libeu.all;
ENTITY LZCounter161Bit IS 
	PORT
	(
		A :  IN  STD_LOGIC_VECTOR(160 DOWNTO 0);
		Z :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END LZCounter161Bit;
ARCHITECTURE Behavioral OF LZCounter161Bit IS 
signal w1499: std_logic;
signal w71: std_logic;
signal w73: std_logic;
signal w33: std_logic;
signal w74: std_logic;
signal w75: std_logic;
signal w34: std_logic;
signal w35: std_logic;
signal w79: std_logic;
signal w1570: std_logic;
signal w1571: std_logic;
signal w1530: std_logic;
signal w1572: std_logic;
signal w1531: std_logic;
signal w1573: std_logic;
signal w1532: std_logic;
signal w1574: std_logic;
signal w1533: std_logic;
signal w1575: std_logic;
signal w1534: std_logic;
signal w1576: std_logic;
signal w1535: std_logic;
signal w1577: std_logic;
signal w1536: std_logic;
signal w1578: std_logic;
signal w1537: std_logic;
signal w1579: std_logic;
signal w1538: std_logic;
signal w1539: std_logic;
signal w1610: std_logic;
signal w1611: std_logic;
signal w1612: std_logic;
signal w1613: std_logic;
signal w1614: std_logic;
signal w1615: std_logic;
signal w1616: std_logic;
signal w1301: std_logic;
signal w1617: std_logic;
signal w1618: std_logic;
signal w1619: std_logic;
signal w1032: std_logic;
signal w1037: std_logic;
signal w481: std_logic;
signal w132: std_logic;
signal w135: std_logic;
signal w1465: std_logic;
signal w40: std_logic;
signal w41: std_logic;
signal w42: std_logic;
signal w45: std_logic;
signal w46: std_logic;
signal w47: std_logic;
signal w216: std_logic;
signal w1580: std_logic;
signal w1581: std_logic;
signal w1540: std_logic;
signal w1582: std_logic;
signal w1500: std_logic;
signal w1541: std_logic;
signal w1501: std_logic;
signal w1583: std_logic;
signal w1542: std_logic;
signal w1584: std_logic;
signal w1502: std_logic;
signal w1543: std_logic;
signal w1503: std_logic;
signal w1585: std_logic;
signal w1544: std_logic;
signal w1586: std_logic;
signal w1545: std_logic;
signal w1504: std_logic;
signal w1505: std_logic;
signal w1587: std_logic;
signal w1546: std_logic;
signal w1588: std_logic;
signal w1547: std_logic;
signal w1506: std_logic;
signal w1507: std_logic;
signal w1233: std_logic;
signal w1589: std_logic;
signal w1548: std_logic;
signal w1549: std_logic;
signal w1508: std_logic;
signal w1509: std_logic;
signal w642: std_logic;
signal w1620: std_logic;
signal w1621: std_logic;
signal w1622: std_logic;
signal w1398: std_logic;
signal w454: std_logic;
signal w100: std_logic;
signal w457: std_logic;
signal w105: std_logic;
signal w147: std_logic;
signal w107: std_logic;
signal w149: std_logic;
signal w109: std_logic;
signal w91: std_logic;
signal w51: std_logic;
signal w10: std_logic;
signal w11: std_logic;
signal w93: std_logic;
signal w14: std_logic;
signal w55: std_logic;
signal w15: std_logic;
signal w16: std_logic;
signal w57: std_logic;
signal w59: std_logic;
signal w846: std_logic;
signal w848: std_logic;
signal w267: std_logic;
signal w1590: std_logic;
signal w1591: std_logic;
signal w1550: std_logic;
signal w1592: std_logic;
signal w1551: std_logic;
signal w1510: std_logic;
signal w1593: std_logic;
signal w1552: std_logic;
signal w1511: std_logic;
signal w1512: std_logic;
signal w1594: std_logic;
signal w1553: std_logic;
signal w1595: std_logic;
signal w1554: std_logic;
signal w1513: std_logic;
signal w1596: std_logic;
signal w1555: std_logic;
signal w1514: std_logic;
signal w1597: std_logic;
signal w1556: std_logic;
signal w1515: std_logic;
signal w1598: std_logic;
signal w1557: std_logic;
signal w1516: std_logic;
signal w1599: std_logic;
signal w1558: std_logic;
signal w1517: std_logic;
signal w1559: std_logic;
signal w1518: std_logic;
signal w1519: std_logic;
signal w1206: std_logic;
signal w1208: std_logic;
signal w615: std_logic;
signal w1010: std_logic;
signal w1054: std_logic;
signal w1056: std_logic;
signal w1059: std_logic;
signal w775: std_logic;
signal w777: std_logic;
signal w110: std_logic;
signal w111: std_logic;
signal w156: std_logic;
signal w116: std_logic;
signal w1482: std_logic;
signal w1444: std_logic;
signal w1487: std_logic;
signal w1176: std_logic;
signal w1135: std_logic;
signal w1139: std_logic;
signal w20: std_logic;
signal w21: std_logic;
signal w22: std_logic;
signal w64: std_logic;
signal w4: std_logic;
signal w25: std_logic;
signal w5: std_logic;
signal w6: std_logic;
signal w69: std_logic;
signal w29: std_logic;
signal w9: std_logic;
signal w272: std_logic;
signal w548: std_logic;
signal w549: std_logic;
signal w277: std_logic;
signal w1560: std_logic;
signal w1561: std_logic;
signal w1520: std_logic;
signal w1562: std_logic;
signal w1521: std_logic;
signal w1563: std_logic;
signal w1522: std_logic;
signal w1564: std_logic;
signal w1523: std_logic;
signal w1565: std_logic;
signal w1524: std_logic;
signal w1566: std_logic;
signal w1525: std_logic;
signal w1567: std_logic;
signal w1526: std_logic;
signal w1568: std_logic;
signal w1527: std_logic;
signal w1569: std_logic;
signal w1528: std_logic;
signal w1529: std_logic;
signal w1299: std_logic;
signal w662: std_logic;
signal w979: std_logic;
signal w668: std_logic;
signal w669: std_logic;
signal w1600: std_logic;
signal w1601: std_logic;
signal w1602: std_logic;
signal w1370: std_logic;
signal w1603: std_logic;
signal w1604: std_logic;
signal w1605: std_logic;
signal w1606: std_logic;
signal w1607: std_logic;
signal w1608: std_logic;
signal w1609: std_logic;
signal w1061: std_logic;
signal w1066: std_logic;
signal w1068: std_logic;
signal w1028: std_logic;
signal w700: std_logic;
signal w470: std_logic;
signal w707: std_logic;
signal w161: std_logic;
signal w120: std_logic;
signal w476: std_logic;
signal w709: std_logic;
signal w122: std_logic;
signal w123: std_logic;
signal w479: std_logic;
signal w124: std_logic;
signal w127: std_logic;
signal w128: std_logic;
signal w129: std_logic;
signal w1451: std_logic;
signal w1492: std_logic;
signal w1411: std_logic;
signal w1413: std_logic;
signal w1495: std_logic;
signal w1414: std_logic;
signal w1496: std_logic;
signal w1456: std_logic;
signal w1497: std_logic;
signal w1457: std_logic;
signal w1498: std_logic;
BEGIN
  w1499 <= w1622 OR w1411;
  w71 <= w1507 OR w59;
  w73 <= w1496 OR w69;
  w33 <= ((w1496 OR (w1496 AND NOT w1595)) OR ((w1496 OR (w1496 AND NOT w1598)) AND NOT w1501)) OR (((w1496 OR (w1496 AND NOT w1569)) OR w979) AND NOT w1497);
  w74 <= w75 AND NOT w1508;
  w75 <= w1496 OR w64;
  w34 <= w35 AND NOT w1503;
  w35 <= ((w1496 OR (w1496 AND NOT w1528)) OR ((w1496 OR (w1496 AND NOT w1531)) AND NOT w1540)) OR (((w1496 OR (w1496 AND NOT w1506)) OR ((w1496 OR w132) AND NOT w1495)) AND NOT w1504);
  w79 <= w1507 AND NOT w1508;
  w1570 <= w1567 OR (A(62) OR A(61));
  w1571 <= w1496 OR w1496;
  w1530 <= w1529 OR (w1527 OR (w1496 OR w1496));
  w1572 <= w1570 OR (w1568 OR (A(58) OR A(57)));
  w1531 <= w1496 OR w1496;
  w1573 <= w1572 OR (w1566 OR (w1565 OR (A(50) OR A(49))));
  w1532 <= w1496 OR w1496;
  w1574 <= A(72) OR A(71);
  w1533 <= w1496 OR w1496;
  w1575 <= A(68) OR A(67);
  w1534 <= w1532 OR (w1496 OR w1496);
  w1576 <= w1574 OR (A(70) OR A(69));
  w1535 <= A(0) OR w1496;
  w1577 <= A(80) OR A(79);
  w1536 <= w1496 OR w1496;
  w1578 <= A(76) OR A(75);
  w1537 <= w1535 OR (w1496 OR w1496);
  w1579 <= w1577 OR (A(78) OR A(77));
  w1538 <= w1537 OR (w1536 OR (w1496 OR w1496));
  w1539 <= w1538 OR (w1534 OR (w1533 OR (w1496 OR w1496)));
  w1610 <= A(144) OR A(143);
  w1611 <= A(140) OR A(139);
  w1612 <= w1610 OR (A(142) OR A(141));
  w1613 <= w1612 OR (w1611 OR (A(138) OR A(137)));
  w1614 <= A(152) OR A(151);
  w1615 <= A(148) OR A(147);
  w1616 <= w1614 OR (A(150) OR A(149));
  w1301 <= (A(136) OR (A(134) AND NOT w1607)) OR ((A(132) OR (A(130) AND NOT w1608)) AND NOT w1609);
  w1617 <= A(160) OR A(159);
  w1618 <= A(156) OR A(155);
  w1619 <= w1617 OR (A(158) OR A(157));
  w1032 <= ((A(80) OR (A(78) AND NOT w1577)) OR ((A(76) OR (A(74) AND NOT w1578)) AND NOT w1579)) OR (((A(72) OR (A(70) AND NOT w1574)) OR ((A(68) OR (A(66) AND NOT w1575)) AND NOT w1576)) AND NOT w1580);
  w1037 <= (w1577 OR (w1578 AND NOT w1579)) OR ((w1574 OR (w1575 AND NOT w1576)) AND NOT w1580);
  w481 <= (w1526 OR (w1527 AND NOT w1529)) OR ((w1521 OR (w1524 AND NOT w1525)) AND NOT w1530);
  w132 <= w1496 AND NOT w1512;
  w135 <= w1508 AND NOT w1513;
  Z(5) <= NOT((w14 OR w15));
  Z(1) <= NOT(w1176);
  w1465 <= (w1587 OR (w1580 AND NOT w1588)) OR ((w1572 OR (w1563 AND NOT w1573)) AND NOT w1589);
  w40 <= w21 OR w22;
  w41 <= w42 AND NOT w1503;
  w42 <= (w1528 OR (w1531 AND NOT w1540)) OR ((w1506 OR (w1512 AND NOT w1495)) AND NOT w1504);
  w45 <= w1501 OR w29;
  w46 <= w47 AND NOT w1503;
  w47 <= w1540 OR (w1495 AND NOT w1504);
  w216 <= (w1496 OR (w1496 AND NOT w1517)) OR ((w1496 OR (w1496 AND NOT w1518)) AND NOT w1519);
  w1580 <= w1579 OR (w1578 OR (A(74) OR A(73)));
  w1581 <= A(88) OR A(87);
  w1540 <= w1528 OR (w1496 OR w1496);
  w1582 <= A(84) OR A(83);
  w1500 <= w1557 OR (w1539 OR w470);
  w1541 <= A(8) OR A(7);
  w1501 <= w1595 OR (w1496 OR w1496);
  w1583 <= w1581 OR (A(86) OR A(85));
  w1542 <= A(4) OR A(3);
  w1584 <= A(96) OR A(95);
  w1502 <= w1569 OR (w1496 OR w1496);
  w1543 <= w1541 OR (A(6) OR A(5));
  w1503 <= w1497 OR (w1502 OR (w1571 OR (w1496 OR w1496)));
  w1585 <= A(92) OR A(91);
  w1544 <= A(16) OR A(15);
  w1586 <= w1584 OR (A(94) OR A(93));
  w1545 <= A(12) OR A(11);
  w1504 <= w1540 OR (w1531 OR (w1496 OR w1496));
  w1505 <= w1496 OR w1496;
  w1587 <= w1586 OR (w1585 OR (A(90) OR A(89)));
  w1546 <= w1544 OR (A(14) OR A(13));
  w1588 <= w1587 OR (w1583 OR (w1582 OR (A(82) OR A(81))));
  w1547 <= w1546 OR (w1545 OR (A(10) OR A(9)));
  w1506 <= w1496 OR w1496;
  w1507 <= w1496 OR w1496;
  w1233 <= (w1593 OR (w1594 AND NOT w1596)) OR ((w1590 OR (w1591 AND NOT w1592)) AND NOT w1597);
  w1589 <= w1588 OR w1028;
  w1548 <= A(24) OR A(23);
  w1549 <= A(20) OR A(19);
  w1508 <= w1505 OR w55;
  w1509 <= w1496 OR w1496;
  w642 <= (w1544 OR (w1545 AND NOT w1546)) OR ((w1541 OR (w1542 AND NOT w1543)) AND NOT w1547);
  w1620 <= w1619 OR (w1618 OR (A(154) OR A(153)));
  w1621 <= w1620 OR (w1616 OR (w1615 OR (A(146) OR A(145))));
  w1622 <= w1621 OR (w1613 OR (w1609 OR (w1608 OR (A(130) OR A(129)))));
  w1398 <= (w1610 OR (w1611 AND NOT w1612)) OR ((w1607 OR (w1608 AND NOT w1609)) AND NOT w1613);
  w454 <= (A(0) OR (w1496 AND NOT w1535)) OR ((w1496 OR (w1496 AND NOT w1536)) AND NOT w1537);
  w100 <= w1496 AND NOT w1510;
  w457 <= (w1496 OR (w1496 AND NOT w1532)) OR ((w1496 OR (w1496 AND NOT w1533)) AND NOT w1534);
  w105 <= w1496 AND NOT w1509;
  w147 <= w1496 OR w1496;
  w107 <= w1510 OR w93;
  w149 <= w1496 OR w1496;
  w109 <= w1496 OR w105;
  Z(6) <= NOT((w1499 OR w20));
  Z(2) <= NOT(((w1456 OR w1457) OR (w1492 AND NOT w1498)));
  w91 <= w1496 OR w1496;
  w51 <= w1504 AND NOT w1503;
  w10 <= w11 AND NOT w1498;
  w11 <= (w1555 OR (w1539 AND NOT w1557)) OR ((w1522 OR (w1503 AND NOT w1523)) AND NOT w1500);
  w93 <= w1496 OR w1496;
  w14 <= w1622 OR (w1589 AND NOT w1499);
  w55 <= w1496 OR w1496;
  w15 <= w16 AND NOT w1498;
  w16 <= w1557 OR (w1523 AND NOT w1500);
  w57 <= w1496 OR w1496;
  w59 <= w1496 OR w1496;
  w846 <= (A(64) OR (A(62) AND NOT w1567)) OR ((A(60) OR (A(58) AND NOT w1568)) AND NOT w1570);
  w848 <= (A(56) OR (A(54) AND NOT w1564)) OR ((A(52) OR (A(50) AND NOT w1565)) AND NOT w1566);
  w267 <= (w216 OR (((w1496 OR w161) OR ((w1496 OR w156) AND NOT w1516)) AND NOT w1520)) OR ((w122 OR w123) AND NOT w1522);
  w1590 <= A(104) OR A(103);
  w1591 <= A(100) OR A(99);
  w1550 <= w1548 OR (A(22) OR A(21));
  w1592 <= w1590 OR (A(102) OR A(101));
  w1551 <= A(32) OR A(31);
  w1510 <= w1496 OR w1496;
  w1593 <= A(112) OR A(111);
  w1552 <= A(28) OR A(27);
  w1511 <= w1509 OR w91;
  w1512 <= w1496 OR w1496;
  w1594 <= A(108) OR A(107);
  w1553 <= w1551 OR (A(30) OR A(29));
  w1595 <= w1496 OR w1496;
  w1554 <= w1553 OR (w1552 OR (A(26) OR A(25)));
  w1513 <= w1511 OR w107;
  w1596 <= w1593 OR (A(110) OR A(109));
  w1555 <= w1554 OR (w1550 OR (w1549 OR (A(18) OR A(17))));
  w1514 <= w1496 OR w1496;
  w1597 <= w1596 OR (w1594 OR (A(106) OR A(105)));
  w1556 <= A(40) OR A(39);
  w1515 <= w1496 OR w1496;
  w1598 <= w1496 OR w1496;
  w1557 <= w1555 OR (w1547 OR (w1543 OR (w1542 OR (A(2) OR A(1)))));
  w1516 <= w1514 OR w147;
  w1599 <= A(120) OR A(119);
  w1558 <= A(36) OR A(35);
  w1517 <= w1496 OR w1496;
  w1559 <= w1556 OR (A(38) OR A(37));
  w1518 <= w1496 OR w1496;
  w1519 <= w1517 OR (w1496 OR w1496);
  w1206 <= (A(128) OR (A(126) AND NOT w1602)) OR ((A(124) OR (A(122) AND NOT w1603)) AND NOT w1604);
  w1208 <= (A(120) OR (A(118) AND NOT w1599)) OR ((A(116) OR (A(114) AND NOT w1600)) AND NOT w1601);
  w615 <= (A(32) OR (A(30) AND NOT w1551)) OR ((A(28) OR (A(26) AND NOT w1552)) AND NOT w1553);
  w1010 <= (A(96) OR (A(94) AND NOT w1584)) OR ((A(92) OR (A(90) AND NOT w1585)) AND NOT w1586);
  w1054 <= (w1010 OR (((A(88) OR (A(86) AND NOT w1581)) OR ((A(84) OR (A(82) AND NOT w1582)) AND NOT w1583)) AND NOT w1587)) OR (w1032 AND NOT w1588);
  w1056 <= (w846 OR (w848 AND NOT w1572)) OR ((w775 OR (w777 AND NOT w1563)) AND NOT w1573);
  w1059 <= ((w1584 OR (w1585 AND NOT w1586)) OR ((w1581 OR (w1582 AND NOT w1583)) AND NOT w1587)) OR (w1037 AND NOT w1588);
  w775 <= (A(48) OR (A(46) AND NOT w1560)) OR ((A(44) OR (A(42) AND NOT w1561)) AND NOT w1562);
  w777 <= (A(40) OR (A(38) AND NOT w1556)) OR ((A(36) OR (A(34) AND NOT w1558)) AND NOT w1559);
  w110 <= w111 AND NOT w1511;
  w111 <= w1496 OR w100;
  w156 <= w1496 AND NOT w1515;
  w116 <= w1510 AND NOT w1511;
  Z(7) <= NOT(w1498);
  Z(3) <= NOT((w4 OR w5));
  w1482 <= (w662 OR (((w454 OR (w457 AND NOT w1538)) OR (w476 AND NOT w1539)) AND NOT w1557)) OR ((w267 OR ((w33 OR w34) AND NOT w1523)) AND NOT w1500);
  w1444 <= w1589 OR (w1573 OR (w1563 OR (w1559 OR (w1558 OR (A(34) OR A(33))))));
  w1487 <= (w668 OR w669) OR ((w272 OR ((w40 OR w41) AND NOT w1523)) AND NOT w1500);
  w1176 <= (w1451 OR ((w1059 OR (w1061 AND NOT w1589)) AND NOT w1499)) OR (w1487 AND NOT w1498);
  w1135 <= (A(112) OR (A(110) AND NOT w1593)) OR ((A(108) OR (A(106) AND NOT w1594)) AND NOT w1596);
  w1139 <= (A(104) OR (A(102) AND NOT w1590)) OR ((A(100) OR (A(98) AND NOT w1591)) AND NOT w1592);
  w20 <= w1500 AND NOT w1498;
  w21 <= w1595 OR (w1598 AND NOT w1501);
  w22 <= w25 AND NOT w1497;
  w64 <= w1496 AND NOT w1507;
  w4 <= ((w1620 OR (w1613 AND NOT w1621)) OR ((w1605 OR (w1597 AND NOT w1606)) AND NOT w1622)) OR (w1465 AND NOT w1499);
  w25 <= w1569 OR (w1571 AND NOT w1502);
  w5 <= w6 AND NOT w1498;
  w6 <= w707 OR (w709 AND NOT w1500);
  w69 <= w1496 AND NOT w1505;
  w29 <= w1502 AND NOT w1497;
  w9 <= (w1621 OR (w1606 AND NOT w1622)) OR ((w1588 OR (w1573 AND NOT w1589)) AND NOT w1499);
  w272 <= ((w1517 OR (w1518 AND NOT w1519)) OR ((w1514 OR (w1515 AND NOT w1516)) AND NOT w1520)) OR ((w127 OR w128) AND NOT w1522);
  w548 <= (A(16) OR (A(14) AND NOT w1544)) OR ((A(12) OR (A(10) AND NOT w1545)) AND NOT w1546);
  w549 <= ((A(8) OR (A(6) AND NOT w1541)) OR ((A(4) OR (A(2) AND NOT w1542)) AND NOT w1543)) AND NOT w1547;
  w277 <= (w1519 OR (w1516 AND NOT w1520)) OR ((w1511 OR w135) AND NOT w1522);
  w1560 <= A(48) OR A(47);
  w1561 <= A(44) OR A(43);
  w1520 <= w1519 OR (w1518 OR (w1496 OR w1496));
  w1562 <= w1560 OR (A(46) OR A(45));
  w1521 <= w1496 OR w1496;
  w1563 <= w1562 OR (w1561 OR (A(42) OR A(41)));
  w1522 <= w1520 OR (w1516 OR (w1515 OR w149));
  w1564 <= A(56) OR A(55);
  w1523 <= w1522 OR (w1513 OR w120);
  w1565 <= A(52) OR A(51);
  w1524 <= w1496 OR w1496;
  w1566 <= w1564 OR (A(54) OR A(53));
  w1525 <= w1521 OR (w1496 OR w1496);
  w1567 <= A(64) OR A(63);
  w1526 <= w1496 OR w1496;
  w1568 <= A(60) OR A(59);
  w1527 <= w1496 OR w1496;
  w1569 <= w1496 OR w1496;
  w1528 <= w1496 OR w1496;
  w1529 <= w1526 OR (w1496 OR w1496);
  w1299 <= (A(144) OR (A(142) AND NOT w1610)) OR ((A(140) OR (A(138) AND NOT w1611)) AND NOT w1612);
  w662 <= (w615 OR (((A(24) OR (A(22) AND NOT w1548)) OR ((A(20) OR (A(18) AND NOT w1549)) AND NOT w1550)) AND NOT w1554)) OR ((w548 OR w549) AND NOT w1555);
  w979 <= (w1496 OR (w1496 AND NOT w1571)) AND NOT w1502;
  w668 <= ((w1551 OR (w1552 AND NOT w1553)) OR ((w1548 OR (w1549 AND NOT w1550)) AND NOT w1554)) OR (w642 AND NOT w1555);
  w669 <= (w479 OR (w481 AND NOT w1539)) AND NOT w1557;
  w1600 <= A(116) OR A(115);
  w1601 <= w1599 OR (A(118) OR A(117));
  w1602 <= A(128) OR A(127);
  w1370 <= (A(160) OR (A(158) AND NOT w1617)) OR ((A(156) OR (A(154) AND NOT w1618)) AND NOT w1619);
  w1603 <= A(124) OR A(123);
  w1604 <= w1602 OR (A(126) OR A(125));
  w1605 <= w1604 OR (w1603 OR (A(122) OR A(121)));
  w1606 <= w1605 OR (w1601 OR (w1600 OR (A(114) OR A(113))));
  w1607 <= A(136) OR A(135);
  w1608 <= A(132) OR A(131);
  w1609 <= w1607 OR (A(134) OR A(133));
  w1061 <= ((w1567 OR (w1568 AND NOT w1570)) OR ((w1564 OR (w1565 AND NOT w1566)) AND NOT w1572)) OR (((w1560 OR (w1561 AND NOT w1562)) OR ((w1556 OR (w1558 AND NOT w1559)) AND NOT w1563)) AND NOT w1573);
  w1066 <= (w1586 OR (w1583 AND NOT w1587)) OR ((w1579 OR (w1576 AND NOT w1580)) AND NOT w1588);
  w1068 <= (w1570 OR (w1566 AND NOT w1572)) OR ((w1562 OR (w1559 AND NOT w1563)) AND NOT w1573);
  w1028 <= w1580 OR (w1576 OR (w1575 OR (A(66) OR A(65))));
  w700 <= ((w1553 OR (w1550 AND NOT w1554)) OR ((w1546 OR (w1543 AND NOT w1547)) AND NOT w1555)) OR (((w1537 OR (w1534 AND NOT w1538)) OR ((w1529 OR (w1525 AND NOT w1530)) AND NOT w1539)) AND NOT w1557);
  w470 <= w1530 OR (w1525 OR (w1524 OR (w1496 OR w1496)));
  w707 <= (w1554 OR (w1547 AND NOT w1555)) OR ((w1538 OR (w1530 AND NOT w1539)) AND NOT w1557);
  w161 <= w1496 AND NOT w1514;
  w120 <= w1508 OR w71;
  w476 <= ((w1496 OR (w1496 AND NOT w1526)) OR ((w1496 OR (w1496 AND NOT w1527)) AND NOT w1529)) OR (((w1496 OR (w1496 AND NOT w1521)) OR ((w1496 OR (w1496 AND NOT w1524)) AND NOT w1525)) AND NOT w1530);
  w709 <= (w1520 OR (w1513 AND NOT w1522)) OR ((w1497 OR w51) AND NOT w1523);
  w122 <= w109 OR w110;
  w123 <= w124 AND NOT w1513;
  w479 <= (w1535 OR (w1536 AND NOT w1537)) OR ((w1532 OR (w1533 AND NOT w1534)) AND NOT w1538);
  w124 <= w73 OR w74;
  w127 <= w1509 OR w116;
  w128 <= w129 AND NOT w1513;
  w129 <= w1505 OR w79;
  Z(4) <= NOT((w9 OR w10));
  Z(0) <= NOT((((w1413 OR w1414) OR ((w1054 OR (w1056 AND NOT w1589)) AND NOT w1499)) OR (w1482 AND NOT w1498)));
  w1451 <= (((w1617 OR (w1618 AND NOT w1619)) OR ((w1614 OR (w1615 AND NOT w1616)) AND NOT w1620)) OR (w1398 AND NOT w1621)) OR ((((w1602 OR (w1603 AND NOT w1604)) OR ((w1599 OR (w1600 AND NOT w1601)) AND NOT w1605)) OR (w1233 AND NOT w1606)) AND NOT w1622);
  w1492 <= w700 OR ((w277 OR ((w45 OR w46) AND NOT w1523)) AND NOT w1500);
  w1411 <= w1606 OR (w1597 OR (w1592 OR (w1591 OR (A(98) OR A(97)))));
  w1413 <= (w1370 OR (((A(152) OR (A(150) AND NOT w1614)) OR ((A(148) OR (A(146) AND NOT w1615)) AND NOT w1616)) AND NOT w1620)) OR ((w1299 OR (w1301 AND NOT w1613)) AND NOT w1621);
  w1495 <= w1506 OR w57;
  w1414 <= ((w1206 OR (w1208 AND NOT w1605)) OR ((w1135 OR (w1139 AND NOT w1597)) AND NOT w1606)) AND NOT w1622;
  w1496 <= '1';
  w1456 <= ((w1619 OR (w1616 AND NOT w1620)) OR ((w1612 OR (w1609 AND NOT w1613)) AND NOT w1621)) OR (((w1604 OR (w1601 AND NOT w1605)) OR ((w1596 OR (w1592 AND NOT w1597)) AND NOT w1606)) AND NOT w1622);
  w1497 <= w1501 OR (w1598 OR (w1496 OR w1496));
  w1457 <= (w1066 OR (w1068 AND NOT w1589)) AND NOT w1499;
  w1498 <= w1499 OR w1444;
END Behavioral;
