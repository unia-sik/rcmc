LIBRARY ieee;
USE ieee.std_logic_1164.all; 
use work.libeu.all;
ENTITY LZCounter53Bit IS 
	PORT
	(
		A :  IN  STD_LOGIC_VECTOR(52 DOWNTO 0);
		Z :  OUT  STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END LZCounter53Bit;
ARCHITECTURE Behavioral OF LZCounter53Bit IS 
signal w21: std_logic;
signal w22: std_logic;
signal w23: std_logic;
signal w26: std_logic;
signal w27: std_logic;
signal w28: std_logic;
signal w321: std_logic;
signal w4: std_logic;
signal w323: std_logic;
signal w5: std_logic;
signal w6: std_logic;
signal w325: std_logic;
signal w326: std_logic;
signal w327: std_logic;
signal w340: std_logic;
signal w328: std_logic;
signal w341: std_logic;
signal w329: std_logic;
signal w342: std_logic;
signal w343: std_logic;
signal w344: std_logic;
signal w345: std_logic;
signal w346: std_logic;
signal w347: std_logic;
signal w348: std_logic;
signal w349: std_logic;
signal w159: std_logic;
signal w174: std_logic;
signal w178: std_logic;
signal w10: std_logic;
signal w198: std_logic;
signal w14: std_logic;
signal w15: std_logic;
signal w16: std_logic;
signal w32: std_logic;
signal w251: std_logic;
signal w253: std_logic;
signal w330: std_logic;
signal w331: std_logic;
signal w332: std_logic;
signal w333: std_logic;
signal w334: std_logic;
signal w335: std_logic;
signal w336: std_logic;
signal w350: std_logic;
signal w337: std_logic;
signal w351: std_logic;
signal w338: std_logic;
signal w339: std_logic;
signal w352: std_logic;
signal w353: std_logic;
signal w354: std_logic;
signal w355: std_logic;
signal w356: std_logic;
signal w181: std_logic;
signal w183: std_logic;
signal w208: std_logic;
BEGIN
  w21 <= w4 OR w5;
  w22 <= w23 AND NOT w330;
  w23 <= (w350 OR (w351 AND NOT w352)) OR ((w333 OR (w339 AND NOT w325)) AND NOT w331);
  w26 <= w328 OR w10;
  w27 <= w28 AND NOT w330;
  w28 <= w352 OR (w325 AND NOT w331);
  w321 <= (A(20) OR (A(18) AND NOT w355)) OR ((A(16) OR (A(14) AND NOT w356)) AND NOT w328);
  w4 <= w355 OR (w356 AND NOT w328);
  w323 <= (A(12) OR (A(10) AND NOT w353)) OR ((A(8) OR (A(6) AND NOT w354)) AND NOT w329);
  w5 <= w6 AND NOT w327;
  w6 <= w353 OR (w354 AND NOT w329);
  w325 <= w333 OR (w326 OR w326);
  w326 <= '1';
  w327 <= w328 OR (w356 OR (A(14) OR A(13)));
  w340 <= w338 OR (w337 OR (A(30) OR A(29)));
  w328 <= w355 OR (A(18) OR A(17));
  Z(0) <= NOT((w198 OR ((w14 OR w15) AND NOT w348)));
  w341 <= A(44) OR A(43);
  w329 <= w353 OR (A(10) OR A(9));
  w342 <= A(40) OR A(39);
  w343 <= w341 OR (A(42) OR A(41));
  w344 <= A(52) OR A(51);
  w345 <= A(48) OR A(47);
  w346 <= w344 OR (A(50) OR A(49));
  w347 <= w346 OR (w345 OR (A(46) OR A(45)));
  Z(2) <= NOT((w208 OR ((w26 OR w27) AND NOT w348)));
  w348 <= w349 OR w174;
  w349 <= w347 OR (w343 OR (w342 OR (A(38) OR A(37))));
  Z(4) <= NOT((w349 OR (w330 AND NOT w348)));
  w159 <= (A(44) OR (A(42) AND NOT w341)) OR ((A(40) OR (A(38) AND NOT w342)) AND NOT w343);
  w174 <= w340 OR (w335 OR (w334 OR (A(22) OR A(21))));
  w178 <= ((A(36) OR (A(34) AND NOT w336)) OR ((A(32) OR (A(30) AND NOT w337)) AND NOT w338)) OR (((A(28) OR (A(26) AND NOT w332)) OR ((A(24) OR (A(22) AND NOT w334)) AND NOT w335)) AND NOT w340);
  w10 <= w329 AND NOT w327;
  w198 <= (((A(52) OR (A(50) AND NOT w344)) OR ((A(48) OR (A(46) AND NOT w345)) AND NOT w346)) OR (w159 AND NOT w347)) OR (w178 AND NOT w349);
  w14 <= w321 OR (w323 AND NOT w327);
  w15 <= w16 AND NOT w330;
  w16 <= w251 OR (w253 AND NOT w331);
  w32 <= w331 AND NOT w330;
  w251 <= (A(4) OR (A(2) AND NOT w350)) OR ((A(0) OR (w326 AND NOT w351)) AND NOT w352);
  w253 <= (w326 OR (w326 AND NOT w333)) OR ((w326 OR (w326 AND NOT w339)) AND NOT w325);
  w330 <= w327 OR (w329 OR (w354 OR (A(6) OR A(5))));
  w331 <= w352 OR (w351 OR (w326 OR w326));
  w332 <= A(28) OR A(27);
  w333 <= w326 OR w326;
  w334 <= A(24) OR A(23);
  w335 <= w332 OR (A(26) OR A(25));
  w336 <= A(36) OR A(35);
  w350 <= A(4) OR A(3);
  w337 <= A(32) OR A(31);
  Z(1) <= NOT(((w181 OR (w183 AND NOT w349)) OR ((w21 OR w22) AND NOT w348)));
  w351 <= A(0) OR w326;
  w338 <= w336 OR (A(34) OR A(33));
  w339 <= w326 OR w326;
  w352 <= w350 OR (A(2) OR A(1));
  w353 <= A(12) OR A(11);
  w354 <= A(8) OR A(7);
  w355 <= A(20) OR A(19);
  w356 <= A(16) OR A(15);
  Z(3) <= NOT(((w347 OR (w340 AND NOT w349)) OR ((w327 OR w32) AND NOT w348)));
  Z(5) <= NOT(w348);
  w181 <= (w344 OR (w345 AND NOT w346)) OR ((w341 OR (w342 AND NOT w343)) AND NOT w347);
  w183 <= (w336 OR (w337 AND NOT w338)) OR ((w332 OR (w334 AND NOT w335)) AND NOT w340);
  w208 <= (w346 OR (w343 AND NOT w347)) OR ((w338 OR (w335 AND NOT w340)) AND NOT w349);
END Behavioral;
