LIBRARY ieee;
USE ieee.std_logic_1164.all; 
use work.libeu.all;
ENTITY LZCounter64Bit IS 
	PORT
	(
		A :  IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		V :  OUT  STD_LOGIC;
		Z :  OUT  STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END LZCounter64Bit;
ARCHITECTURE Behavioral OF LZCounter64Bit IS 
signal w21: std_logic;
signal w24: std_logic;
signal w25: std_logic;
signal w26: std_logic;
signal w2: std_logic;
signal w320: std_logic;
signal w3: std_logic;
signal w4: std_logic;
signal w322: std_logic;
signal w323: std_logic;
signal w324: std_logic;
signal w325: std_logic;
signal w326: std_logic;
signal w8: std_logic;
signal w88: std_logic;
signal w327: std_logic;
signal w340: std_logic;
signal w328: std_logic;
signal w341: std_logic;
signal w342: std_logic;
signal w329: std_logic;
signal w343: std_logic;
signal w344: std_logic;
signal w345: std_logic;
signal w346: std_logic;
signal w347: std_logic;
signal w348: std_logic;
signal w349: std_logic;
signal w157: std_logic;
signal w174: std_logic;
signal w12: std_logic;
signal w197: std_logic;
signal w14: std_logic;
signal w15: std_logic;
signal w16: std_logic;
signal w30: std_logic;
signal w250: std_logic;
signal w19: std_logic;
signal w34: std_logic;
signal w330: std_logic;
signal w318: std_logic;
signal w331: std_logic;
signal w332: std_logic;
signal w333: std_logic;
signal w334: std_logic;
signal w335: std_logic;
signal w336: std_logic;
signal w350: std_logic;
signal w337: std_logic;
signal w351: std_logic;
signal w338: std_logic;
signal w352: std_logic;
signal w339: std_logic;
signal w147: std_logic;
signal w180: std_logic;
signal w182: std_logic;
signal w207: std_logic;
signal w20: std_logic;
BEGIN
  w21 <= (w346 OR (w347 AND NOT w348)) OR ((w329 OR (w332 AND NOT w322)) AND NOT w327);
  w24 <= w324 OR w8;
  w25 <= w26 AND NOT w326;
  w26 <= w348 OR (w322 AND NOT w327);
  w2 <= w351 OR (w352 AND NOT w324);
  w320 <= (A(23) OR (A(21) AND NOT w349)) OR ((A(19) OR (A(17) AND NOT w350)) AND NOT w325);
  w3 <= w4 AND NOT w323;
  w4 <= w349 OR (w350 AND NOT w325);
  w322 <= w329 OR (A(5) OR A(4));
  w323 <= w324 OR (w352 OR (A(25) OR A(24)));
  w324 <= w351 OR (A(29) OR A(28));
  w325 <= w349 OR (A(21) OR A(20));
  w326 <= w323 OR (w325 OR (w350 OR (A(17) OR A(16))));
  w8 <= w325 AND NOT w323;
  w88 <= (A(39) OR (A(37) AND NOT w328)) OR ((A(35) OR (A(33) AND NOT w330)) AND NOT w331);
  w327 <= w348 OR (w347 OR (A(9) OR A(8)));
  w340 <= A(63) OR A(62);
  w328 <= A(39) OR A(38);
  Z(0) <= NOT((w197 OR ((w14 OR w15) AND NOT w344)));
  w341 <= A(59) OR A(58);
  w342 <= w340 OR (A(61) OR A(60));
  w329 <= A(7) OR A(6);
  w343 <= w342 OR (w341 OR (A(57) OR A(56)));
  w344 <= w345 OR (w336 OR (w331 OR (w330 OR (A(33) OR A(32)))));
  w345 <= w343 OR (w339 OR (w338 OR (A(49) OR A(48))));
  w346 <= A(15) OR A(14);
  w347 <= A(11) OR A(10);
  Z(2) <= NOT((w207 OR ((w24 OR w25) AND NOT w344)));
  w348 <= w346 OR (A(13) OR A(12));
  w349 <= A(23) OR A(22);
  Z(4) <= NOT((w345 OR (w326 AND NOT w344)));
  w157 <= (A(55) OR (A(53) AND NOT w337)) OR ((A(51) OR (A(49) AND NOT w338)) AND NOT w339);
  w174 <= ((A(63) OR (A(61) AND NOT w340)) OR ((A(59) OR (A(57) AND NOT w341)) AND NOT w342)) OR (w157 AND NOT w343);
  w12 <= w327 OR (w322 OR (w332 OR (A(1) OR A(0))));
  w197 <= w174 OR ((((A(47) OR (A(45) AND NOT w333)) OR ((A(43) OR (A(41) AND NOT w334)) AND NOT w335)) OR (w88 AND NOT w336)) AND NOT w345);
  w14 <= w318 OR (w320 AND NOT w323);
  w15 <= w16 AND NOT w326;
  w16 <= w250 OR (((A(7) OR (A(5) AND NOT w329)) OR w147) AND NOT w327);
  w30 <= w327 AND NOT w326;
  w250 <= (A(15) OR (A(13) AND NOT w346)) OR ((A(11) OR (A(9) AND NOT w347)) AND NOT w348);
  w19 <= w2 OR w3;
  w34 <= A(37) OR A(36);
  V <= NOT((w344 OR (w326 OR w12)));
  w330 <= A(35) OR A(34);
  w318 <= (A(31) OR (A(29) AND NOT w351)) OR ((A(27) OR (A(25) AND NOT w352)) AND NOT w324);
  w331 <= w328 OR w34;
  w332 <= A(3) OR A(2);
  w333 <= A(47) OR A(46);
  w334 <= A(43) OR A(42);
  w335 <= w333 OR (A(45) OR A(44));
  w336 <= w335 OR (w334 OR (A(41) OR A(40)));
  w350 <= A(19) OR A(18);
  w337 <= A(55) OR A(54);
  Z(1) <= NOT(((w180 OR (w182 AND NOT w345)) OR ((w19 OR w20) AND NOT w344)));
  w351 <= A(31) OR A(30);
  w338 <= A(51) OR A(50);
  w352 <= A(27) OR A(26);
  w339 <= w337 OR (A(53) OR A(52));
  Z(3) <= NOT(((w343 OR (w336 AND NOT w345)) OR ((w323 OR w30) AND NOT w344)));
  w147 <= (A(3) OR (A(1) AND NOT w332)) AND NOT w322;
  Z(5) <= NOT(w344);
  w180 <= (w340 OR (w341 AND NOT w342)) OR ((w337 OR (w338 AND NOT w339)) AND NOT w343);
  w182 <= (w333 OR (w334 AND NOT w335)) OR ((w328 OR (w330 AND NOT w331)) AND NOT w336);
  w207 <= (w342 OR (w339 AND NOT w343)) OR ((w335 OR (w331 AND NOT w336)) AND NOT w345);
  w20 <= w21 AND NOT w326;
END Behavioral;
